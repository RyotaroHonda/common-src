library ieee;
use ieee.std_logic_1164.all;

package defMiiRstTimer is
  constant kWidthPhyAddr  : positive:= 5;

  constant kWidthCounter  : positive:= 28;

end package defMiiRstTimer;

